module multi-clock()

endmodule 